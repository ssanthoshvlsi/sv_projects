class generator;
    transaction tr;
    mailbox #(transaction) mbxgd;

