module axi_slave(
        input clk,
        input resetn,
        //write address channel
        input awvalid,//master send new address
        output reg awready,//slave is ready to accept request
        input [3:0] awid, //unique id for txn
        input [3:0] awlen, //burst length 1 to 16 //burst length = awlenth + 1 beats   
        input [2:0] awsize, //2^awsize //1,2,4,8,16,...128 unique transaction size
        input [31:0] awaddr,//write addr
        input [1:0] awburst,//burst type fixed, incr, wrap//000, 001, 010
        //write data channel
        input wvalid,//master sending to slave newdata
        output reg wready,//slave is ready to accept new data
        input [3:0] wid,//unique id for fpr txns
        input [31:0] wdata,//data
        input [3:0] wstrb,//lane having valid data
        input wlast,//last trnx in write data
        //write reponse 
        input bready,
        output reg bvalid,
        output reg [3:0] bid,
        output reg [1:0] bresp,
        //read address channel
        output reg arready,
        input [3:0] arid,
        input [31:0] araddr,
        input [3:0] arlen,
        input [2:0] arsize,
        input [1:0] arburst,
        input arvalid,
        //read data channel
        output reg [3:0] rid,
        output reg [31:0] rdata,
        output reg [1:0] rresp,
        output reg rlast,
        output reg rvalid,
        input rready
);
typedef enum bit[1:0]{awidle = 2'b00, awstart = 2'b01, awready = 2'b10} awstate_type;
awstate_type awstate, awnext_state;
reg[31:0] awaddrt;
//reset decoder
always_ff @(posedge clk, negedge resetn) begin
        if(!resetn) begin
                awstate <= awidle;//write addr fsm
                wstart <= widle;//write data fsm
                bstate <= bidle;//write response
        end
        else begin
                awstate <= awnext_state;
                wstate <= wnext_state;
                bstate <= bnext_state;
        end
end
//fsm for write address channel
always_comb begin
        case(awstate)
                awidle: begin
                        awready = 1'b0;
                        awnext_state = awstart;
                end
                awstart: begin
                        if(awvalid) begin
                                awnext_state = awready;
                                awaddrt = awaddr;
                        end
                        else 
                                awnext_state = awstart;
                end
                awready: begin
                        awready = 1'b1;
                        awnext_state = awidle;
                end
        endcase
end
//fsm for write data channel
reg [31:0] wdatat;
reg [7:0] mem[128] = '{default:12};
reg [31:0] retaddr;
reg [31:0] nextaddr;
reg first;
//compute next addr during fixed
function bit[31:0] data_wr_fixed(input[3:0] wstrb, input[31:0] awaddrt);
        unique case(wstrb)
        4'b0001 : begin
                mem[awaddrt] = wdatat[7:0];
        end
        4'b0010 : begin
                mem[awaddrt] = wdatat[15:8];
        end
        4'b0011 : begin 
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[15:8];
        end
        4'b0100 : begin
                mem[awaddrt] = wdatat[23:16];
        end
        4'b0101 : begin 
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[23:16];
        end
        4'b0110 : begin 
                mem[awaddrt] = wdatat[15:8];
                mem[awaddrt + 1] = wdatat[23:16];
        end
        4'b0111 : begin 
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[15:8];
                mem[awaddrt + 2] = wdatat[23:16];
        end
        4'b1000 : begin
                mem[awaddrt] = wdatat[31:24];
        end
        4'b1001 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[31:24];
        end
        4'b1010 : begin
                mem[awaddrt] = wdatat[15:8];
                mem[awaddrt + 1] = wdatat[31:24];
        end
        4'b1011 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[15:8];
                mem[awaddrt + 2] = wdatat[31:24];
        end
        4'b1100 : begin
                mem[awaddrt] = wdatat[23:16];
                mem[awaddrt + 1] = wdatat[31:24];
        end
        4'b1101 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[23:16];
                mem[awaddrt + 2] = wdatat[31:24];
        end
        4'b1110 : begin
                mem[awaddrt] = wdatat[15:0];
                mem[awaddrt + 1] = wdatat[23:16];
                mem[awaddrt + 2] = wdatat[31:24];
        end
        4'b1111 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[15:8];
                mem[awaddrt + 2] = wdatat[23:16];
                mem[awaddrt + 3] = wdatat[31:24];
        end
endcase
return awaddrt;
endfunction
//compute address during INCR burst type
function bit[31:0] data_wr_incr(input[3:0] wstrb, input[31:0] awaddrt);
        bit[31:0] addr;
        unique case(wstrb)
        4'b0001 : begin
                mem[awaddrt] = wdatat[7:0];
                addr = awaddrt + 1;
        end
        4'b0010 : begin
                mem[awaddrt] = wdatat[15:8];
                addr = awaddrt + 1;
        end
        4'b0011 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[15:8];
                addr = awaddrt + 2;
        end
        4'b0100 : begin
                mem[awaddrt] = wdatat[23:16];
                addr = awaddrt + 1;
        end
        4'b0101 : begin 
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[23:16];
                addr = awaddrt + 2;
        end
        4'b0110 : begin 
                mem[awaddrt] = wdatat[15:8];
                mem[awaddrt + 1] = wdatat[23:16];
                addr = awaddrt + 2;
        end
        4'b0111 : begin 
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[15:8];
                mem[awaddrt + 2] = wdatat[23:16];
                addr = awaddrt + 3;
        end
        4'b1000 : begin
                mem[awaddrt] = wdatat[31:24];
                addr = awaddrt + 1;
        end
        4'b1001 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[31:24];
                addr = awaddrt + 2;
        end
        4'b1010 : begin
                mem[awaddrt] = wdatat[15:8];
                mem[awaddrt + 1] = wdatat[31:24];
                addr = awaddrt + 2;
        end
        4'b1011 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[15:8];
                mem[awaddrt + 2] = wdatat[31:24];
                addr = awaddrt + 3;
        end
        4'b1100 : begin
                mem[awaddrt] = wdatat[23:16];
                mem[awaddrt + 1] = wdatat[31:24];
                addr = awaddrt + 2;
        end
        4'b1101 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[23:16];
                mem[awaddrt + 2] = wdatat[31:24];
                addr = awaddrt + 3;
        end
        4'b1110 : begin
                mem[awaddrt] = wdatat[15:0];
                mem[awaddrt + 1] = wdatat[23:16];
                mem[awaddrt + 2] = wdatat[31:24];
                addr = awaddrt + 3;
        end
        4'b1111 : begin
                mem[awaddrt] = wdatat[7:0];
                mem[awaddrt + 1] = wdatat[15:8];
                mem[awaddrt + 2] = wdatat[23:16];
                mem[awaddrt + 3] = wdatat[31:24];
                addr = awaddrt + 4;
        end
endcase
return awaddrt;
endfunction
//compute WRAP boundary
function bit[7:0] wrap_boundary(input bit[3:0] awlen, input bit[2:0] awsize);
        bit[7:0] boundary;
        unique case(awlen)
        4'b0001 : begin
                unique case(awsize)
                3'b000 : begin
                        boundary = 2 * 1;
                end
                3'b001 : begin
                        boundary = 2 * 2;
                end
                3'b010 : begin
                        boundary = 2 * 4;
                end
                endcase
        end
        4'b0011 : begin
                unique case(awsize)
                3'b000 : begin
                        boundary = 4 * 1;
                end
                3'b001 : begin
                        boundary = 4 * 2;
                end
                3'b010 : begin
                        boundary = 4 * 4;
                end
                endcase
        end
        4'b0111 : begin
                unique case(awsize)
                3'b000 : begin
                        boundary = 8 * 1;
                end
                3'b001 : begin
                        boundary = 8 * 2;
                end
                3'b010 : begin
                        boundary = 8 * 4;
                end
                endcase
        end
        4'b1111 : begin
                unique case(awsize)
                3'b000 : begin
                        boundary = 16 * 1;
                end
                3'b001 : begin
                        boundary = 16 * 2;
                end
                3'b010 : begin
                        boundary = 16 * 4;
                end
                endcase
        end
        endcase
        return boundary;
endfunction
function bit[31:0] data_wr_wrap(input[3:0] wstrb, input[31:0] awaddrt, input[7:0] wboundary);
    bit[31:0] addr1, addr2, addr3, addr4;
    bit[31:0] nextaddr, nextaddr2;
    unique case(wstrb)
    4'b0001 : begin
             mem[awaddrt] = wdatat[7:0];
             if((awaddrt + 1) % wboundary == 0)
                 addr1 = (awaddrt + 1) - wboundary;
             else
                 addr1 = awaddrt + 1;
    return addr1;
    end
    4'b0010 : begin
            mem[awaddrt] = wdatat[15:8];
            if((awaddrt + 1) % wboundary == 0)
               addr1 = (awaddrt + 1) - wboundary;
            else
               addr1 = awaddrt + 1;
    return addr1;
    end
    4'b0011 : begin
            mem[awaddrt] = wdatat[7:0];
            if((awaddrt + 1) % wboundary == 0)
               addr1 = (awaddrt + 1) - wboundary;
            else
               addr1 = awaddrt + 1;
            mem[addr1] = wdatat[15:8];
            if(addr1 + 1) % wboundary == 0)
              addr2 = (addr1 + 1) - wboundary;
            else
              addr2 = addr1 + 1;
    return addr2; 
    end
    4'b0100 : begin
            mem[awaddrt] = wdatat[23:16];
            if((awaddrt + 1) % wboundary == 0)
             addr1 = (awaddrt + 1) - wboundary;
            else
             addr1 = awaddrt + 1;
   return addr1;
   end
   4'b0101 : begin 
           mem[awaddrt] = wdatat[7:0];
            if((awaddrt + 1) % wboundary == 0)
               addr1 = (awaddrt + 1) - wboundary;
            else
               addr1 = awaddrt + 1;
           mem[addr1] = wdatat[23:16];
             if(addr1 + 1) % wboundary == 0)
              addr2 = (addr1 + 1) - wboundary;
              else
              addr2 = addr1 + 1;
   return addr2; 
   end
   4'b0110 : begin 
           mem[awaddrt] = wdatat[15:8];
            if((awaddrt + 1) % wboundary == 0)
               addr1 = (awaddrt + 1) - wboundary;
            else
               addr1 = awaddrt + 1;
           mem[addr1] = wdatat[23:16];
            if(addr1 + 1) % wboundary == 0)
              addr2 = (addr1 + 1) - wboundary;
            else
              addr2 = addr1 + 1;
   return addr2; 
   end
   4'b0111 : begin 
           mem[awaddrt] = wdatat[7:0];
           if((awaddrt + 1) % wboundary == 0)
            addr1 = (awaddrt + 1) - wboundary;
           else
            addr1 = awaddrt + 1;
           mem[addr1] = wdatat[15:8];
           if((addr1 + 1) % wboundary == 0)
            addr2 = (addr1 + 1) - wboundary;
           else
            addr2 = addr1 + 1;
           mem[addr2] = wdatat[23:16];
           if((addr2 + 1) % wboundary == 0)
            addr3 = (addr2 + 1) - wboundary;
           else
            addr3 = addr2 + 1;
   return addr3;
   end
   4'b1000 : begin
           mem[awaddrt] = wdatat[31:24];
           if((awaddrt + 1) % wboundary == 0)
           addr1 = (awaddrt + 1) - wboundary;
           else
           addr1 = awaddrt + 1;
   return addr1;
   end
   4'b1001 : begin
           mem[awaddrt] = wdatat[7:0];
           if((awaddrt + 1) % wboundary == 0)
            addr1 = (awaddrt + 1) - wboundary;
           else
           addr1 = awaddrt + 1;
           mem[addr1] = wdatat[31:24];
           if((addr1 + 1) % wboundary == 0)
            addr2 = (addr1 + 1) - wboundary;
           else
            addr2 = addr1 + 1;
   return addr2;
   end
   4'b1010 : begin
           mem[awaddrt] = wdatat[15:8];
           if((awaddrt + 1) % wboundary == 0)
            addr1 = (awaddrt + 1) - wboundary;
           else
           addr1 = awaddrt + 1;
           mem[addr1] = wdatat[31:24];
           if((addr1 + 1) % wboundary == 0)
            addr2 = (addr1 + 1) - wboundary;
           else
            addr2 = addr1 + 1;
   return addr2;
   end
   4'b1011 : begin
           mem[awaddrt] = wdatat[7:0];
           if((awaddrt + 1) % wboundary == 0)
            addr1 = (awaddrt + 1) - wboundary;
           else
           addr1 = awaddrt + 1;
           mem[addr1] = wdatat[15:8];
           if((addr1 + 1) % wboundary == 0)
            addr2 = (addr1 + 1) - wboundary;
           else
            addr2 = addr1 + 1;
           mem[addr2] = wdatat[31:24];
           if((addr2 + 1) % wboundary == 0)
            addr3 = (addr2 + 1) - wboundary;
           else
            addr3 = addr2 + 1;
   return addr3;
   end
   4'b1100 : begin
           mem[awaddrt] = wdatat[23:16];
           if((awaddrt + 1) % wboundary == 0)
            addr1 = (awaddrt + 1) - wboundary;
           else
           addr1 = awaddrt + 1;
           mem[addr1] = wdatat[31:24];
           if((addr1 + 1) % wboundary == 0)
            addr2 = (addr1 + 1) - wboundary;
           else
            addr2 = addr1 + 1;
   return addr2;
   end
   4'b1101 : begin
           mem[awaddrt] = wdatat[7:0];
           if((awaddrt + 1) % wboundary == 0)
            addr1 = (awaddrt + 1) - wboundary;
           else
           addr1 = awaddrt + 1;
           mem[addr1] = wdatat[23:16];
           if((addr1 + 1) % wboundary == 0)
            addr2 = (addr1 + 1) - wboundary;
           else
            addr2 = addr1 + 1;
           mem[addr2] = wdatat[31:24];
           if((addr2 + 1) % wboundary == 0)
            addr3 = (addr2 + 1) - wboundary;
           else
            addr3 = addr2 + 1;
   return addr3;
   end
   4'b1110 : begin
           mem[awaddrt] = wdatat[15:0];
           if((awaddrt + 1) % wboundary == 0)
            addr1 = (awaddrt + 1) - wboundary;
           else
           addr1 = awaddrt + 1;
           mem[addr1] = wdatat[23:16];
           if((addr1 + 1) % wboundary == 0)
            addr2 = (addr1 + 1) - wboundary;
           else
            addr2 = addr1 + 1;
           mem[addr2] = wdatat[31:24];
           if((addr2 + 1) % wboundary == 0)
            addr3 = (addr2 + 1) - wboundary;
           else
            addr3 = addr2 + 1;
   return addr3;
   end
   4'b1111 : begin
           mem[awaddrt] = wdatat[7:0];
           if((awaddrt + 1) % wboundary == 0)
            addr1 = (awaddrt + 1) - wboundary;
           else
           addr1 = awaddrt + 1;
           mem[addr1] = wdatat[15:8];
           if((addr1 + 1) % wboundary == 0)
            addr2 = (addr1 + 1) - wboundary;
           else
            addr2 = addr1 + 1;
           mem[addr2] = wdatat[23:16];
           if((addr2 + 1) % wboundary == 0)
            addr3 = (addr2 + 1) - wboundary;
           else
            addr3 = addr2 + 1;
           mem[addr3] = wdatat[31:24];
           if((addr3 + 1) % wboundary == 0)
            addr4 = (addr3 + 1) - wboundary;
           else
            addr4 = addr3 + 1;
   return addr4;
   end
endcase
endfunction
reg[7:0] boundary;
reg[3:0] wlen_count;
typedef enum bit[2:0]{widle = 0, wstart = 1, wready = 2, wvalid = 3, waddr_dec = 4} wstate_type;
wstate_type wstate, wnext_state;
always_comb begin
    case(wstate)
        widle: begin
            wready = 1'b0;
            wnext_state = wstart;
            first = 1'b0;
            wlen_count = 0;
        end
        wstart: begin
            if(wvalid) begin
                wnext_state = waddr_dec;
                wdatat = wdata;
            end
            else begin
                wnext_state = wstart;
            end
        end
        waddr_dec: begin
            wnext_state = wready;
            if(first == 0) begin
                nextaddr = awaddr;
                first = 1'b1;
            end
            else if(wlen_count != (awlen + 1)) begin
                nextaddr = retaddr;
            end
            else begin
                nextaddr = awaddr;
            end
        end
        wready: begin
            if(wlast == 1'b1) begin
                wnext_state = widle;
                wready = 1'b0;
                wlen_count = 0;
                first = 0;
            end
            else begin
                wnext_state = wvalid;
                wready = 1'b1;
            end
            case(awburst)
                2'b00: begin//fixed mode
                    retaddr = data_wr_fixed(wstrb, awaddr);
                end
                2'b01: begin//inc mode
                    retaddr = data_wr_incr(wstrb, nextaddr);
                end
                2'b10: begin//wrap mode
                    boundary = wrap_boundary(awlen, awsize);//calculating wrapping boundary
                    retaddr = data_wr_wrap(wstrb, nextaddr, boundary);//generate next address
                end
            endcase
        end
        wvalid: begin
            wready = 1'b0;
            wnext_state = wstart;
            if(wlen_count != (awlen + 1))
                wlen_count = wlen_count + 1;
            else 
                wlen_count = wlen_count;
        end
    endcase
end
    //fsm for write response
typedef enum bit[1:0]{bidle = 0, bdetect_last = 1, bstart = 2, bwait = 3} bstate_type;
bstate_type bstart, bnext_state;
always_comb begin
    case(bstate)
        bidle: begin
            bid = 1'b0;
            bresp = 1'b0;
            bvalid = 1'b0;
            bnext_state = bdetect_last;
        end
        bdetect_last: begin
            if(wlast)
                bnext_state = bstart;
            else
                bnext_state = bdetect_last;
        end
        bstart: begin
            bid = awid;
            bvalid = 1'b1;
            bnext_state = bwait;
            if((awaddr < 128) && (awsize <= 3'b011))
                bresp = 2'b00;//okay
            else if(awsize > 3'b011)
                bresp = 2'b10;//slverr
            else
                bresp = 2'b11;//no slave addr
        end
        bwait: begin
            if(bready == 1'b1)
                bnext_state = bidle;
            else 
                bnext_state = bwait;
        end
    endcase
end
//fsm read address
//read data in fixed mode
function void read_data_fixed(input [31:0]addr, input[2:0] arsize);
    unique case(arsize)
    3'b000: begin
        rdata[7:0] = mem[addr];
    end
    3'b001: begin
        rdata[7:0] = mem[addr];
        rdata[15:8] = mem[addr + 1];
    end
    3'b010: begin
        rdata[7:0] = mem[addr];
        rdata[15:8] = mem[addr + 1];
        rdata[23:16] = mem[addr + 2];
        rdata[31:24] = mem[addr + 3];
    end
    endcase
endfunction
//read data in incr mode
function bit[31:0] read_data_incr(input [31:0] addr, input[2:0] arsize);
    bit[31:0] nextaddr;
    unique case(arsize)
    3'b000: begin
        rdata[7:0] = mem[addr];
        nextaddr = addr + 1;
    end
    3'b001: begin
        rdata[7:0] = mem[addr];
        rdata[15:8] = mem[addr + 1];
        nextaddr = addr + 2;
    end
    3'b010: begin
        rdata[7:0] = mem[addr];
        rdata[15:8] = mem[addr + 1];
        rdata[23:16] = mem[addr + 2];
        nextaddr = addr + 3;
    end






endmodule
interface axi_if();
        //write address channel
        logic awvalid;//master send new address
        logic awready;//slave is ready to accept request
        logic [3:0] awid; //unique id for txn
        logic [3:0] awlen; //burst length 1 to 16 //burst length = awlenth + 1 beats   
        logic [2:0] awsize; //2^awsize //1;2;4;8;16;...128 unique transaction size
        logic [31:0] awaddr;//write addr
        logic [1:0] awburst;//burst type fixed; incr; wrap//000; 001; 010
        //write data channel
        logic wvalid;//master sending to slave newdata
        logic wready;//slave is ready to accept new data
        logic [3:0] wid;//unique id for fpr txns
        logic [31:0] wdata;//data
        logic [3:0] wstrb;//lane having valid data
        logic wlast;//last trnx in write data
        //write reponse 
        logic bready;
        logic bvalid;
        logic [3:0] bid;
        logic [1:0] bresp;
        //read address channel
        logic arready;
        logic [3:0] arid;
        logic [31:0] araddr;
        logic [3:0] arlen;
        logic [2:0] arsize;
        logic [1:0] arburst;
        logic arvalid;
        //read data channel
        logic [3:0] rid;
        logic [31:0] rdata;
        logic [1:0] rresp;
        logic rlast;
        logic rvalid;
        logic rready;
        logic clk;
        logic resetn;
        logic [31:0] addr_wrapwr;
        logic [31:0] addr_wraprd;
endinterface
